//---------------------------------------------------------------------- 
// File Name: sk_buff_pkg.svh
// Author: dzplay
// Email: dzplay@qq.com
// Date: 2023.09.28
// MD5: 8d45881764a4ed4e17c03743f2cea131
//---------------------------------------------------------------------- 
`ifndef SKBUFF_PKG_SV
`define SKBUFF_PKG_SV

package libs_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "skbuff.sv"

endpackage

`endif