//---------------------------------------------------------------------- 
// File Name: libs_pkg.svh
// Author: dzplay
// Email: dzplay@qq.com
// Date: 2024.07.16
// MD5: 8d45881764a4ef2cea131d4e17c03743
//---------------------------------------------------------------------- 

`ifndef LIBS_PKG_SV
`define LIBS_PKG_SV

package libs_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "libs.sv"

endpackage

`endif
