//---------------------------------------------------------------------- 
// File Name: wheels_pkg.svh
// Author: dzplay
// Email: dzplay@qq.com
// Date: 2024.07.16
// MD5: 8d45881764a4ef2cea131d4e17c03743
//---------------------------------------------------------------------- 

`ifndef WHEELS_PKG_SV
`define WHEELS_PKG_SV

package wheels_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "wheels.sv"

endpackage

`endif
