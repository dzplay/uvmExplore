// filelist version 1.0
// -------------------------------------------------------------
// $SIM_ROOT/common/avalon_module/src/burst_read_master.v
// +incdir+$SIM_ROOT/common/avalon_module/verif/avalon_agent
// $SIM_ROOT/common/avalon_module/verif/avalon_agent/avalon_if.sv
// $SIM_ROOT/common/avalon_module/verif/avalon_agent/avalon_pkg.svh
// +incdir+$SIM_ROOT/common/avalon_module/verif/env
// $SIM_ROOT/common/avalon_module/verif/env/tb_env_pkg.svh
// +incdir+$SIM_ROOT/common/avalon_module/verif/tests
// $SIM_ROOT/common/avalon_module/verif/tests/test_base.sv
// +incdir+$SIM_ROOT/common/avalon_module/verif
// $SIM_ROOT/common/avalon_module/verif/tb_top.sv
// -fsdb
// -------------------------------------------------------------
// filelist version 2.0
// -------------------------------------------------------------
// -f $SIM_ROOT/common/avalon_module/verif/tb_top.f
// -fsdb
// -------------------------------------------------------------

`undef EXPLICIT_MON
// `include "tb_top.sv"
