//---------------------------------------------------------------------- 
// File Name: pcap_pkg.svh
// Author: dzplay
// Email: dzplay@qq.com
// Date: 2023.09.28
// MD5: 8d45881764a4ed4e17c03743f2cea131
//---------------------------------------------------------------------- 
`ifndef PCAP_PKG_SV
`define PCAP_PKG_SV

package libs_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "pcap.sv"

endpackage

`endif